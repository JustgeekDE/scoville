*** Simple full adder ***

* Supply
Vs VCC GND dc 5V ac 0V

* First XOR
QXA1 VCC XA1b XA1e BC547B
QXA2 XA1e XA2b XA2e BC547B
QXA3 XA3c XA3b GND BC547B
QXA4 XA3c XA4b GND BC547B
QXA5 XA5c XA5b GND BC547B
QXA6 XA5c XA6b GND BC547B

RXA1 B XA1b 10k
RXA2 INV XA2b 10k
RXA3 B XA3b 10k
RXA4 INV XA4b 10k
RXA5 XA2e XA5b 10k
RXA6 XA3c XA6b 10k
RXA7 XA2e GND 10k
RXA8 VCC XA3c 10k
RXA9 VCC XA5c 1k

* Second XOR
QXB1 VCC XB1b XB1e BC547B
QXB2 XB1e XB2b XB2e BC547B
QXB3 XB3c XB3b GND BC547B
QXB4 XB3c XB4b GND BC547B
QXB5 XOR XB5b GND BC547B
QXB6 XOR XB6b GND BC547B

RXB1 A XB1b 10k
RXB2 XA5c XB2b 10k
RXB3 A XB3b 10k
RXB4 XA5c XB4b 10k
RXB5 XB2e XB5b 10k
RXB6 XB3c XB6b 10k
RXB7 XB2e GND 10k
RXB8 VCC XB3c 10k
RXB9 VCC XOR 1k

* Third XOR
QXC1 VCC XC1b XC1e BC547B
QXC2 XC1e XC2b XC2e BC547B
QXC3 XC3c XC3b GND BC547B
QXC4 XC3c XC4b GND BC547B
QXC5 CARRY XC5b GND BC547B
QXC6 CARRY XC6b GND BC547B

RXC1 XOR XC1b 10k
RXC2 C XC2b 10k
RXC3 XOR XC3b 10k
RXC4 C XC4b 10k
RXC5 XC2e XC5b 10k
RXC6 XC3c XC6b 10k
RXC7 XC2e GND 10k
RXC8 VCC XC3c 10k
RXC9 VCC CARRY 1k

* NAND
QNA1 NAND NA1b GND BC547B
RNA1 XB2e NA1b 10k
RNA2 VCC NAND 1k

* OR
QOA1 OA1c OA1b GND BC547B
QOA2 OA1c OA2b GND BC547B
QOA3 SUM OA3b GND BC547B

ROA1 XB2e OA1b 10k
ROA2 XC2e OA2b 10k
ROA3 OA1c OA3b 10k
ROA4 VCC OA1c 10k
ROA5 VCC SUM 10k


.model BC547B NPN ()

.end
