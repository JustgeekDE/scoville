*** Basic ALU ***
Q1 VCC N002 N007 BC547B
Q2 N007 N010 AND_X1 BC547B
R1 AND_X1 GND 1k
R2 VCC NOR_X1 1k
R3 N002 B 10K
R4 N010 INV 10k
R5 N019 B 10k
R6 N022 INV 10k
R7 N013 AND_X1 10k
R8 N016 NOR_X1 10k
R9 VCC XOR_X1 1k
Q3 NOR_X1 N019 GND BC547B
Q4 NOR_X1 N022 GND BC547B
Q5 XOR_X1 N013 GND BC547B
Q6 XOR_X1 N016 GND BC547B
Q7 VCC N003 N008 BC547B
Q8 N008 N011 AND_X2 BC547B
R10 AND_X2 GND 1k
R11 VCC NOR 1k
R12 N003 A 10K
R13 N011 XOR_X1 10k
R14 N020 A 10k
R15 N023 XOR_X1 10k
R16 N014 AND_X2 10k
R17 N017 NOR 10k
R18 VCC XOR 1k
Q9 NOR N020 GND BC547B
Q10 NOR N023 GND BC547B
Q11 XOR N014 GND BC547B
Q12 XOR N017 GND BC547B
Q13 VCC N004 N009 BC547B
Q14 N009 N012 AND_X3 BC547B
R19 AND_X3 GND 1k
R20 VCC NOR_X3 1k
R21 N004 XOR 10K
R22 N012 C 10k
R23 N021 XOR 10k
R24 N024 C 10k
R25 N015 AND_X3 10k
R26 N018 NOR_X3 10k
R27 VCC SUM 1k
Q15 NOR_X3 N021 GND BC547B
Q16 NOR_X3 N024 GND BC547B
Q17 SUM N015 GND BC547B
Q18 SUM N018 GND BC547B
R28 VCC N005 1k
Q19 N005 AND_X2 GND BC547B
Q20 N005 AND_X3 GND BC547B
R29 N006 N005 10K
Q21 CARRY N006 GND BC547B
R30 VCC CARRY 1k
R31 N001 AND_X2 10K
Q22 NAND N001 GND BC547B
R32 VCC NAND 1k

Vs VCC GND dc 5V ac 0V
.model BC547B NPN ()

.end
