*** Simple NAND ***

* Supply
Vs VCC GND dc 5V ac 0V

* Transistors
Qa out aBase aEm BC547B
Ra inA aBase 10k

Qb aBase bBase GND BC547B
Rb inB bBase 10k

* Pullup
Rpull VCC out 10k

.model BC547B NPN ()

.end
