*** Basic XOR ***

* Supply
Vs VCC GND dc 5V ac 0V

* AND
QA1 VCC A1b A1e BC547B
QA2 A1e A2b AND BC547B

RA1 A A1b 10k
RA2 B A2b 10k
RA3 AND GND 1k

* FIRST NOR
QB1 NOR B1b GND BC547B
QB2 NOR B2b GND BC547B

RB1 VCC NOR 1k
RB2 A B1b 10k
RB3 B B2b 10k

* SECOND NOR
QC1 XOR C1b GND BC547B
QC2 XOR C2b GND BC547B

RC1 VCC XOR 1k
RC2 AND C1b 10k
RC3 NOR C2b 10k

.model BC547B NPN ()

.end
